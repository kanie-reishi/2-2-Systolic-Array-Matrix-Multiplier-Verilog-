library verilog;
use verilog.vl_types.all;
entity tb_systolic_2x2 is
end tb_systolic_2x2;
